// 100 MHz scale
`timescale 10ns/10ns

module top_tb;
endmodule
