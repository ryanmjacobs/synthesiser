module clkdiv_tb;
endmodule
